
module FastFourierTransform( 
//clk, reset
//									  input [:0] s0,input [:0] s1, input [:0] s2, input [:0] s3, input [:0] s4, input [:0] s4, input [:0] s5, input [:0] s6, input [:0] s7, input [:0] s8, input [:0] s9,
//									  input [:0] s10, input [:0] s11, input [:0] s12, input [:0] s13, input [:0] s14, input [:0] s15, output [:0] x0, output [:0] x1, output [:0] x2 , output [:0] x3, 
//									  output [:0] x4, output [:0] x5, output [:0] x6, output [:0] x7, output [:0] x8 , output [:0] x9, output [:0] x10, output [:0] x11, output [:0] x12, output [:0] x13,
//									  output [:0] x14, output [:0] x15, output [:0] x16

);
//	// ASSIGN THE TWIDDLE FACTORs
//	assign W0 =
//	assign W1 = 
//	assign W2 = 
//	assign W3 =
//	assign W4 = 
//	assign w5 = 
//	assign w6 =
//	assign w7 =
//	
//	enum logic [2:0] {halt, stage1, stage2, stage3, stage4 } curr_state, next_state;
//	
//	logic [:0]  butterflyinput0 ,butterflyinput1, butterflyinput2, butterflyinput3, butterflyinput4, butterflyinput5, butterflyinput6, butterflyinput7;
//
//	always_ff@(posedge clk or posedge reset)
//		begin
//			if (reset)
//				curr_state = halt
//			else 
//				
//				
//		
//		
//		
//		end
//		
//		
//		
//		
endmodule 